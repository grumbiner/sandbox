netcdf VIIRS_winds {
//---------
dimensions:
//---------
	BufferSize = 36158 ;
	SizeOne = 1 ;

//---------
variables:
//---------

// This is the first array

	int Time(BufferSize) ;
		Time:long_name = "date/time of measurement" ;
		Time:coordinates = "Time Latitude Longitude Altitude" ;
		Time:units = "secs since 1970-01-01 00:00:00" ;
		Time:_FillValue = -999 ;
	float Latitude(BufferSize) ;
		Latitude:long_name = "Wind Latitude" ;
		Latitude:coordinates = "Time Latitude Longitude Altitude" ;
		Latitude:units = "degrees_north" ;
		Latitude:_FillValue = -999.f ;
		Latitude:valid_range = -90.f, 90.f ;
	float Longitude(BufferSize) ;
		Longitude:long_name = "Wind Longitude" ;
		Longitude:coordinates = "Time Latitude Longitude Altitude" ;
		Longitude:units = "degrees_east" ;
		Longitude:_FillValue = -999.f ;
		Longitude:valid_range = -180.f, 180.f ;
	float Wind_Speed(BufferSize) ;
		Wind_Speed:long_name = "Speed of average wind vector (m/s)" ;
		Wind_Speed:coordinates = "Time Latitude Longitude Altitude" ;
		Wind_Speed:units = "m.s-1" ;
		Wind_Speed:_FillValue = -999.f ;
		Wind_Speed:valid_range = 0.f, 155.f ;
	float Wind_Dir(BufferSize) ;
		Wind_Dir:long_name = "Direction of average wind vector (degrees)" ;
		Wind_Dir:coordinates = "Time Latitude Longitude Altitude" ;
		Wind_Dir:units = "degree" ;
		Wind_Dir:_FillValue = -999.f ;
		Wind_Dir:valid_range = 0.f, 360.f ;
	float UComponent1(BufferSize) ;
		UComponent1:long_name = "u-component of first (reverse time) vector" ;
		UComponent1:coordinates = "Time Latitude Longitude Altitude" ;
		UComponent1:units = "m.s-1" ;
		UComponent1:_FillValue = -999.f ;
	float VComponent1(BufferSize) ;
		VComponent1:long_name = "v-component of first (reverse time) vector" ;
		VComponent1:coordinates = "Time Latitude Longitude Altitude" ;
		VComponent1:units = "m.s-1" ;
		VComponent1:_FillValue = -999.f ;
	float UComponent2(BufferSize) ;
		UComponent2:long_name = "u-component of second (forward) vector" ;
		UComponent2:coordinates = "Time Latitude Longitude Altitude" ;
		UComponent2:units = "m.s-1" ;
		UComponent2:_FillValue = -999.f ;
	float VComponent2(BufferSize) ;
		VComponent2:long_name = "v-component of second (forward) vector" ;
		VComponent2:coordinates = "Time Latitude Longitude Altitude" ;
		VComponent2:units = "m.s-1" ;
		VComponent2:_FillValue = -999.f ;
	float MedianPress(BufferSize) ;
		MedianPress:long_name = "Pressure assignment of tracer (mb)" ;
		MedianPress:coordinates = "Time Latitude Longitude Altitude" ;
		MedianPress:units = "hPa" ;
		MedianPress:_FillValue = -999.f ;
		MedianPress:valid_range = 0.f, 1100.f ;
	float Altitude(BufferSize) ;
		Altitude:long_name = "Derived altitude of tracer from pressure (m)" ;
		Altitude:coordinates = "Time Latitude Longitude Altitude" ;
		Altitude:units = "m" ;
		Altitude:_FillValue = -999.f ;
		Altitude:valid_range = -300.f, 30000.f ;
	float Fcst_Spd(BufferSize) ;
		Fcst_Spd:long_name = "speed of forecast" ;
		Fcst_Spd:coordinates = "Time Latitude Longitude Altitude" ;
		Fcst_Spd:units = "m.s-1" ;
		Fcst_Spd:_FillValue = -999.f ;
	float Fcst_Dir(BufferSize) ;
		Fcst_Dir:long_name = "direction of forecast" ;
		Fcst_Dir:coordinates = "Time Latitude Longitude Altitude" ;
		Fcst_Dir:units = "degree" ;
		Fcst_Dir:_FillValue = -999.f ;
	float CorrCoeff(BufferSize) ;
		CorrCoeff:long_name = "Correlation coefficient of first vector" ;
		CorrCoeff:coordinates = "Time Latitude Longitude Altitude" ;
		CorrCoeff:units = "1" ;
		CorrCoeff:_FillValue = -999.f ;
	float CorrCoeff2(BufferSize) ;
		CorrCoeff2:long_name = "Correlation coefficient of second vector" ;
		CorrCoeff2:coordinates = "Time Latitude Longitude Altitude" ;
		CorrCoeff2:units = "1" ;
		CorrCoeff2:_FillValue = -999.f ;
	float MedianBT(BufferSize) ;
		MedianBT:long_name = "Representative BrtTemp of tracer" ;
		MedianBT:coordinates = "Time Latitude Longitude Altitude" ;
		MedianBT:units = "Kelvin" ;
		MedianBT:_FillValue = -999.f ;
	float ExpectedErr(BufferSize) ;
		ExpectedErr:long_name = "Expected Error" ;
		ExpectedErr:coordinates = "Time Latitude Longitude Altitude" ;
		ExpectedErr:units = "m.s-1" ;
		ExpectedErr:_FillValue = -999.f ;
	int QI(BufferSize) ;
		QI:long_name = "Quality Indicator (QI) of derived wind (0-100, with 100 being the best)" ;
		QI:coordinates = "Time Latitude Longitude Altitude" ;
		QI:units = "1" ;
		QI:_FillValue = -98 ;
		QI:valid_range = 1, 100 ;
	int QISpdFlag(BufferSize) ;
		QISpdFlag:long_name = "QI test - Speed Consistency Flag" ;
		QISpdFlag:coordinates = "Time Latitude Longitude Altitude" ;
		QISpdFlag:units = "1" ;
		QISpdFlag:_FillValue = -999 ;
	int QIDirFlag(BufferSize) ;
		QIDirFlag:long_name = "QI test - Direction Consistency Flag" ;
		QIDirFlag:coordinates = "Time Latitude Longitude Altitude" ;
		QIDirFlag:units = "1" ;
		QIDirFlag:_FillValue = -999 ;
	int QIVecFlag(BufferSize) ;
		QIVecFlag:long_name = "QI test - Vector Consistency Flag" ;
		QIVecFlag:coordinates = "Time Latitude Longitude Altitude" ;
		QIVecFlag:units = "1" ;
		QIVecFlag:_FillValue = -999 ;
	int QILocConsistencyFlg(BufferSize) ;
		QILocConsistencyFlg:long_name = "QI test - Buddy Consistency(cloest neighbor) Flag" ;
		QILocConsistencyFlg:coordinates = "Time Latitude Longitude Altitude" ;
		QILocConsistencyFlg:units = "1" ;
		QILocConsistencyFlg:_FillValue = -999 ;
	int QIFcstFlag(BufferSize) ;
		QIFcstFlag:long_name = "QI test - Forecast Consistency Flag" ;
		QIFcstFlag:coordinates = "Time Latitude Longitude Altitude" ;
		QIFcstFlag:units = "1" ;
		QIFcstFlag:_FillValue = -999 ;
	float VariancePress(BufferSize) ;
		VariancePress:long_name = "Standard deviation of cloud top pressure values in target scene (hPa)" ;
		VariancePress:coordinates = "Time Latitude Longitude Altitude" ;
		VariancePress:units = "hPa" ;
		VariancePress:_FillValue = -999.f ;
	float SatZen(BufferSize) ;
		SatZen:long_name = "satellite zenith angle" ;
		SatZen:coordinates = "Time Latitude Longitude Altitude" ;
		SatZen:units = "degree" ;
		SatZen:_FillValue = -999.f ;
	float LatMatch(BufferSize) ;
		LatMatch:long_name = "Latitude of the match in the preceding image" ;
		LatMatch:coordinates = "Time Latitude Longitude Altitude" ;
		LatMatch:units = "degrees_north" ;
		LatMatch:_FillValue = -999.f ;
	float LonMatch(BufferSize) ;
		LonMatch:long_name = "Longitude of the match in the preceding image" ;
		LonMatch:coordinates = "Time Latitude Longitude Altitude" ;
		LonMatch:units = "degrees_east" ;
		LonMatch:_FillValue = -999.f ;
	float LatMatch2(BufferSize) ;
		LatMatch2:long_name = "Latitude of the match in the succeeding image" ;
		LatMatch2:coordinates = "Time Latitude Longitude Altitude" ;
		LatMatch2:units = "degrees_north" ;
		LatMatch2:_FillValue = -999.f ;
	float LonMatch2(BufferSize) ;
		LonMatch2:long_name = "Longitude of the match in the succeeding image" ;
		LonMatch2:coordinates = "Time Latitude Longitude Altitude" ;
		LonMatch2:units = "degrees_east" ;
		LonMatch2:_FillValue = -999.f ;
	int PointIndex(BufferSize) ;
		PointIndex:long_name = "Cold sample counter in brightness temperature histogram" ;
		PointIndex:coordinates = "Time Latitude Longitude Altitude" ;
		PointIndex:units = "1" ;
		PointIndex:_FillValue = -999 ;
	float StdDevMVD1(BufferSize) ;
		StdDevMVD1:long_name = "Standard deviation of largest 5x5 cluster (sample 1 - reverse vector)" ;
		StdDevMVD1:coordinates = "Time Latitude Longitude Altitude" ;
		StdDevMVD1:units = "1" ;
		StdDevMVD1:_FillValue = -999.f ;
	float StdDevMVD2(BufferSize) ;
		StdDevMVD2:long_name = "Standard deviation of largest 5x5 cluster (sample 2 - forward vector)" ;
		StdDevMVD2:coordinates = "Time Latitude Longitude Altitude" ;
		StdDevMVD2:units = "1" ;
		StdDevMVD2:_FillValue = -999.f ;
	float PctOfAvg1(BufferSize) ;
		PctOfAvg1:long_name = "Standard deviation of sample 1 divided by magnitude of average displacement" ;
		PctOfAvg1:coordinates = "Time Latitude Longitude Altitude" ;
		PctOfAvg1:units = "1" ;
		PctOfAvg1:_FillValue = -999.f ;
	float PctOfAvg2(BufferSize) ;
		PctOfAvg2:long_name = "Standard deviation of sample 2 divided by magnitude of average displacement" ;
		PctOfAvg2:coordinates = "Time Latitude Longitude Altitude" ;
		PctOfAvg2:units = "1" ;
		PctOfAvg2:_FillValue = -999.f ;
	int NumClusters1(BufferSize) ;
		NumClusters1:long_name = "Number of distinct motion clusters from DBSCAN analysis  (sample 1 - reverse vector)" ;
		NumClusters1:coordinates = "Time Latitude Longitude Altitude" ;
		NumClusters1:units = "1" ;
		NumClusters1:_FillValue = -999 ;
	int NumClusters2(BufferSize) ;
		NumClusters2:long_name = "Number of distinct motion clusters from DBSCAN analysis  (sample 2 - forward vector)" ;
		NumClusters2:coordinates = "Time Latitude Longitude Altitude" ;
		NumClusters2:units = "1" ;
		NumClusters2:_FillValue = -999 ;
	int MaxClusterSize1(BufferSize) ;
		MaxClusterSize1:long_name = "Size of largest DBSCAN cluster (sample 1 - reverse vector)" ;
		MaxClusterSize1:coordinates = "Time Latitude Longitude Altitude" ;
		MaxClusterSize1:units = "1" ;
		MaxClusterSize1:_FillValue = -999 ;
	int MaxClusterSize2(BufferSize) ;
		MaxClusterSize2:long_name = "Size of largest DBSCAN cluster (sample 2 - forward vector)" ;
		MaxClusterSize2:coordinates = "Time Latitude Longitude Altitude" ;
		MaxClusterSize2:units = "1" ;
		MaxClusterSize2:_FillValue = -999 ;
	int LandFlag(BufferSize) ;
		LandFlag:long_name = "Land Mask" ;
		LandFlag:coordinates = "Time Latitude Longitude Altitude" ;
		LandFlag:units = "1" ;
		LandFlag:_FillValue = -999 ;
	int InversionFlag(BufferSize) ;
		InversionFlag:long_name = "Low-level inversion flag" ;
		InversionFlag:coordinates = "Time Latitude Longitude Altitude" ;
		InversionFlag:units = "1" ;
		InversionFlag:_FillValue = -999 ;
	int CloudPhase(BufferSize) ;
		CloudPhase:long_name = "Dominant cloud phase of target scene" ;
		CloudPhase:coordinates = "Time Latitude Longitude Altitude" ;
		CloudPhase:units = "1" ;
		CloudPhase:_FillValue = -999 ;
	int CloudType(BufferSize) ;
		CloudType:long_name = "Dominant cloud type of target scene" ;
		CloudType:coordinates = "Time Latitude Longitude Altitude" ;
		CloudType:units = "1" ;
		CloudType:_FillValue = -999 ;
	float TempGrad(BufferSize) ;
		TempGrad:long_name = "NWP vertical temperature gradient (+/- 200 hPa about pressure assignment of tracer)" ;
		TempGrad:coordinates = "Time Latitude Longitude Altitude" ;
		TempGrad:units = "Kelvin" ;
		TempGrad:_FillValue = -999.f ;
	float Wind_Speed_Shear(BufferSize) ;
		Wind_Speed_Shear:long_name = "NWP vertical wind shear (+/- 200 hPa about pressure assignment of tracer)" ;
		Wind_Speed_Shear:coordinates = "Time Latitude Longitude Altitude" ;
		Wind_Speed_Shear:units = "m.s-1" ;
		Wind_Speed_Shear:_FillValue = -999.f ;
	float MinCTP(BufferSize) ;
		MinCTP:long_name = "Minimum cloud-top pressure (hPa) in largest cluster" ;
		MinCTP:coordinates = "Time Latitude Longitude Altitude" ;
		MinCTP:units = "hPa" ;
		MinCTP:_FillValue = -999.f ;
	float MaxCTP(BufferSize) ;
		MaxCTP:long_name = "Maximum cloud-top pressure (hPa) in largest cluster" ;
		MaxCTP:coordinates = "Time Latitude Longitude Altitude" ;
		MaxCTP:units = "hPa" ;
		MaxCTP:_FillValue = -999.f ;
	float MinCTT(BufferSize) ;
		MinCTT:long_name = "Minimum cloud-top temperature (K) in largest cluster" ;
		MinCTT:coordinates = "Time Latitude Longitude Altitude" ;
		MinCTT:units = "Kelvin" ;
		MinCTT:_FillValue = -999.f ;
	float MaxCTT(BufferSize) ;
		MaxCTT:long_name = "Maximum cloud-top temperature (K) in largest cluster" ;
		MaxCTT:coordinates = "Time Latitude Longitude Altitude" ;
		MaxCTT:units = "Kelvin" ;
		MaxCTT:_FillValue = -999.f ;
	float CombinedMedianHgtErr(BufferSize) ;
		CombinedMedianHgtErr:long_name = "Representative height error (hPa)" ;
		CombinedMedianHgtErr:coordinates = "Time Latitude Longitude Altitude" ;
		CombinedMedianHgtErr:units = "hPa" ;
		CombinedMedianHgtErr:_FillValue = -999.f ;
	float CombinedMedianTempErr(BufferSize) ;
		CombinedMedianTempErr:long_name = "Representative temperature error" ;
		CombinedMedianTempErr:coordinates = "Time Latitude Longitude Altitude" ;
		CombinedMedianTempErr:units = "Kelvin" ;
		CombinedMedianTempErr:_FillValue = -999.f ;
	int Flag(BufferSize) ;
		Flag:long_name = "Internal Quality Flag" ;
		Flag:coordinates = "Time Latitude Longitude Altitude" ;
		Flag:units = "1" ;
		Flag:_FillValue = -99 ;
		Flag:valid_range = 0, 16 ;
	int PriorImageDate(BufferSize) ;
		PriorImageDate:long_name = "Date(Year+Julian day) of prior image" ;
		PriorImageDate:coordinates = "" ;
		PriorImageDate:units = "1" ;
		PriorImageDate:_FillValue = 0 ;
	int PriorImageTime(BufferSize) ;
		PriorImageTime:long_name = "Time(HHMM) of prior image" ;
		PriorImageTime:coordinates = "" ;
		PriorImageTime:units = "1" ;
		PriorImageTime:_FillValue = 0 ;
	int NextImageDate(BufferSize) ;
		NextImageDate:long_name = "Date(Year+Julian day) of subsequent image" ;
		NextImageDate:coordinates = "" ;
		NextImageDate:units = "1" ;
		NextImageDate:_FillValue = 0 ;
	int NextImageTime(BufferSize) ;
		NextImageTime:long_name = "Time(HHMM) of subsequent image" ;
		NextImageTime:coordinates = "" ;
		NextImageTime:units = "1" ;
		NextImageTime:_FillValue = 0 ;
	int NumTargets_Total(SizeOne);
		NumTargets_Total:long_name = "Total targets identified" ;
		NumTargets_Total:units = "1" ;
	int SatID(SizeOne) ;
		SatID:long_name = "Satellite ID" ;
		SatID:units = "1" ;
	int AMVChannel(SizeOne) ;
		AMVChannel:long_name = "Channel number" ;
		AMVChannel:units = "1" ;
	int TimeInterval(SizeOne) ;
		TimeInterval:long_name = "minutes between images" ;
		TimeInterval:units = "1" ;
	int BoxSize(SizeOne) ;
		BoxSize:long_name = "Target box size being tracked" ;
		BoxSize:units = "1" ;
	int LagSize(SizeOne) ;
		LagSize:long_name = "Lag size(in pixels)" ;
		LagSize:units = "1" ;
	int NestedTrackingFlg(SizeOne) ;
		NestedTrackingFlg:long_name = "Nested tracking flag" ;
		NestedTrackingFlg:units = "1" ;
	int Target_Type(SizeOne) ;
		Target_Type:long_name = "Target type(0=clear; 1=cloudy)" ;
		Target_Type:units = "1" ;
	int NumOfChn(SizeOne) ;
		NumOfChn:long_name = "Number of Channels" ;
		NumOfChn:units = "1" ;
	int NumQAVals(SizeOne) ;
		NumQAVals:long_name = "Number of QA Flag Values" ;
		NumQAVals:units = "1" ;
	float QA_Value_0(SizeOne) ;
		QA_Value_0:long_name = "% of QA flag value of 0: good wind; passes all QC checks" ;
		QA_Value_0:units = "1" ;
	float QA_Value_1(SizeOne) ;
		QA_Value_1:long_name = "% of QA flag value of 1: Maximum gradient below acceptable threshold" ;
		QA_Value_1:units = "1" ;
	float QA_Value_2(SizeOne) ;
		QA_Value_2:long_name = "% of QA flag value of 2: Target located on earth edge" ;
		QA_Value_2:units = "1" ;
	float QA_Value_3(SizeOne) ;
		QA_Value_3:long_name = "% of QA flag value of 3: Cloud amount failures(less than 10% cloud cover for cloud track winds or greater than 0% cloud cover for water vapor clear sky winds)" ;
		QA_Value_3:units = "1" ;
	float QA_Value_4(SizeOne) ;
		QA_Value_4:long_name = "% of QA flag value of 4: Median pressure not found" ;
		QA_Value_4:units = "1" ;
	float QA_Value_5(SizeOne) ;
		QA_Value_5:long_name = "% of QA flag value of 5: Bad or missing brightness temperature in target scene" ;
		QA_Value_5:units = "1" ;
	float QA_Value_6(SizeOne) ;
		QA_Value_6:long_name = "% of QA flag value of 6: More than 1 cloud layer present" ;
		QA_Value_6:units = "1" ;
	float QA_Value_7(SizeOne) ;
		QA_Value_7:long_name = "% of QA flag value of 7: Target scene too coherent (not enough structure for reliable tracking)" ;
		QA_Value_7:units = "1" ;
	float QA_Value_8(SizeOne) ;
		QA_Value_8:long_name = "% of QA flag value of 8: Tracking correlation below 0.6 (not used for nested tracking)" ;
		QA_Value_8:units = "1" ;
	float QA_Value_9(SizeOne) ;
		QA_Value_9:long_name = "% of QA flag value of 9: u-component acceleration greater than 5 m/s (for winds generated from visible channel) or 10 m/s (for winds generated from any other channel)" ;
		QA_Value_9:units = "1" ;
	float QA_Value_10(SizeOne) ;
		QA_Value_10:long_name = "% of QA flag value of 10: v-component acceleration greater than 5 m/s (for winds generated from visible channel) or 10 m/s (for winds generated from any other channel)" ;
		QA_Value_10:units = "1" ;
	float QA_Value_11(SizeOne) ;
		QA_Value_11:long_name = "% of QA flag value of 11: u- and v- component accelerations greater than 5 m/s (for winds generated from visible channel) or 10 m/s (for winds generated from any other channel)" ;
		QA_Value_11:units = "1" ;
	float QA_Value_12(SizeOne) ;
		QA_Value_12:long_name = "% of QA flag value of 12: Derived wind slower than 3 m/s" ;
		QA_Value_12:units = "1" ;
	float QA_Value_13(SizeOne) ;
		QA_Value_13:long_name = "% of QA flag value of 13: Target scene too close to day/night terminator (visible and SWIR only)" ;
		QA_Value_13:units = "1" ;
	float QA_Value_14(SizeOne) ;
		QA_Value_14:long_name = "% of QA flag value of 14: Median pressure used for height assignment outside acceptable pressure range (channel dependent)" ;
		QA_Value_14:units = "1" ;
	float QA_Value_15(SizeOne) ;
		QA_Value_15:long_name = "% of QA flag value of 15: Match found on boundary of search region" ;
		QA_Value_15:units = "1" ;
	float QA_Value_16(SizeOne) ;
		QA_Value_16:long_name = "% of QA flag value of 16: Gross difference from forecast wind (channel dependent)" ;
		QA_Value_16:units = "1" ;
	float QA_Value_17(SizeOne) ;
		QA_Value_17:long_name = "% of QA flag value of 17: Median pressure of largest cluster for first image pair is too different from median pressure of largest cluster for second image pair  only valid for nested tracking" ;
		QA_Value_17:units = "1" ;
	float QA_Value_18(SizeOne) ;
		QA_Value_18:long_name = "% of QA flag value of 18: Search region extends beyond domain of data buffer" ;
		QA_Value_18:units = "1" ;
	float QA_Value_19(SizeOne) ;
		QA_Value_19:long_name = "% of QA flag value of 19: Expected Error (EE) too high" ;
		QA_Value_19:units = "1" ;
	float QA_Value_20(SizeOne) ;
		QA_Value_20:long_name = "% of QA flag value of 20: Missing data in search box" ;
		QA_Value_20:units = "1" ;
	float QA_Value_21(SizeOne) ;
		QA_Value_21:long_name = "% of QA flag value of 21: No winds are available for the clustering algorithm" ;
		QA_Value_21:units = "1" ;
	float QA_Value_22(SizeOne) ;
		QA_Value_22:long_name = "% of QA flag value of 22: No clusters were found" ;
		QA_Value_22:units = "1" ;
	float WndSpdMean(SizeOne) ;
		WndSpdMean:long_name = "Mean of target wind speed" ;
		WndSpdMean:units = "m/s" ;
	float WndSpdMin(SizeOne) ;
		WndSpdMin:long_name = "Min of target wind speed" ;
		WndSpdMin:units = "m.s-1" ;
	float WndSpdMax(SizeOne) ;
		WndSpdMax:long_name = "Max of target wind speed" ;
		WndSpdMax:units = "m.s-1" ;
	float WndSpdStdDev(SizeOne) ;
		WndSpdStdDev:long_name = "StdDev of target wind speed" ;
		WndSpdStdDev:units = "m.s-1" ;
	int NumOfAtmosLayers(SizeOne) ;
		NumOfAtmosLayers:long_name = "Number of atmospheric layers" ;
		NumOfAtmosLayers:units = "1" ;
	int NumGoodWnds_Layer1(SizeOne) ;
		NumGoodWnds_Layer1:long_name = "Number of good winds for atmospheric layer1(100 - 399.9 mb)" ;
		NumGoodWnds_Layer1:units = "1" ;
	int NumGoodWnds_Layer2(SizeOne) ;
		NumGoodWnds_Layer2:long_name = "Number of good winds for atmospheric layer2(400 - 699.9 mb)" ;
		NumGoodWnds_Layer2:units = "1" ;
	int NumGoodWnds_Layer3(SizeOne) ;
		NumGoodWnds_Layer3:long_name = "Number of good winds for atmospheric layer3(700 - 1000 mb)" ;
		NumGoodWnds_Layer3:units = "1" ;
	float CldHgtMean_Layer1(SizeOne) ;
		CldHgtMean_Layer1:long_name = "cloud height mean for atmospheric layer1" ;
		CldHgtMean_Layer1:units = "hPa" ;
	float CldHgtMean_Layer2(SizeOne) ;
		CldHgtMean_Layer2:long_name = "cloud height mean for atmospheric layer2" ;
		CldHgtMean_Layer2:units = "hPa" ;
	float CldHgtMean_Layer3(SizeOne) ;
		CldHgtMean_Layer3:long_name = "cloud height mean for atmospheric layer3" ;
		CldHgtMean_Layer3:units = "hPa" ;
	float CldHgtMin_Layer1(SizeOne) ;
		CldHgtMin_Layer1:long_name = "cloud height min for atmospheric layer1" ;
		CldHgtMin_Layer1:units = "hPa" ;
	float CldHgtMin_Layer2(SizeOne) ;
		CldHgtMin_Layer2:long_name = "cloud height min for atmospheric layer2" ;
		CldHgtMin_Layer2:units = "hPa" ;
	float CldHgtMin_Layer3(SizeOne) ;
		CldHgtMin_Layer3:long_name = "cloud height min for atmospheric layer3" ;
		CldHgtMin_Layer3:units = "hPa" ;
	float CldHgtMax_Layer1(SizeOne) ;
		CldHgtMax_Layer1:long_name = "cloud height max for atmospheric layer1" ;
		CldHgtMax_Layer1:units = "hPa" ;
	float CldHgtMax_Layer2(SizeOne) ;
		CldHgtMax_Layer2:long_name = "cloud height max for atmospheric layer2" ;
		CldHgtMax_Layer2:units = "hPa" ;
	float CldHgtMax_Layer3(SizeOne) ;
		CldHgtMax_Layer3:long_name = "cloud height max for atmospheric layer3" ;
		CldHgtMax_Layer3:units = "hPa" ;
	float CldHgtStdDev_Layer1(SizeOne) ;
		CldHgtStdDev_Layer1:long_name = "Standard deviation about mean height (hPa) assigned to good derived winds in atmospheric layer 1" ;
		CldHgtStdDev_Layer1:units = "hPa" ;
	float CldHgtStdDev_Layer2(SizeOne) ;
		CldHgtStdDev_Layer2:long_name = "Standard deviation about mean height (hPa) assigned to good derived winds in atmospheric layer 2" ;
		CldHgtStdDev_Layer2:units = "hPa" ;
	float CldHgtStdDev_Layer3(SizeOne) ;
		CldHgtStdDev_Layer3:long_name = "Standard deviation about mean height (hPa) assigned to good derived winds in atmospheric layer 3" ;
		CldHgtStdDev_Layer3:units = "hPa" ;
	float WndSpdStdDev_Layer1(SizeOne) ;
		WndSpdStdDev_Layer1:long_name = "Standard deviation about mean wind speed (m/s) assigned to good derived winds in atmospheric layer 1" ;
		WndSpdStdDev_Layer1:units = "m.s-1" ;
	float WndSpdStdDev_Layer2(SizeOne) ;
		WndSpdStdDev_Layer2:long_name = "Standard deviation about mean wind speed (m/s) assigned to good derived winds in atmospheric layer 2" ;
		WndSpdStdDev_Layer2:units = "m.s-1" ;
	float WndSpdStdDev_Layer3(SizeOne) ;
		WndSpdStdDev_Layer3:long_name = "Standard deviation about mean wind speed (m/s) assigned to good derived winds in atmospheric layer 3" ;
		WndSpdStdDev_Layer3:units = "m.s-1" ;

// This is the last array

	float GoodWndClrCld(SizeOne) ;
		GoodWndClrCld:long_name = "% of good winds for Clear/Cloudy sky" ;
		GoodWndClrCld:units = "1" ;

//------------------
// global attributes:
//------------------
		:Title = "AWG_NOP_AMV" ;
		:Source = "AIT_Framework" ;
}
