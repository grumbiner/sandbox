//----------------------------------------------------------------------------
//
// QSS Group
//
//
// NAME:
//       aot_geo.cdl
//
// PURPOSE:
//       netCDF4 file specification for VIIRS MOD GEO file.
//
//       This file specification document is written in the network Common
//       Data Form Language (CDL) to define NetCDF dimension names and
//       sizes, and to declare attributes and arrays in terms of the
//       dimensions.
//
// CATEGORY:
//       VIIRS: Data Storage
//
// LANGUAGE:
//       CDL
//
// RESTRICTIONS:
//       None
//
// EXAMPLE:
//       This file specification should be used with the ncgen utility to
//       produce the initial (empty) file for VIIRS granule data:
//
//           $ ncgen -b -k3 aot_geo.cdl
//
//
// MODIFICATION HISTORY:
//       Written by:   Yi Song, IMSG, 12/29/09
//                     Yi.Song@noaa.gov
//
//  $Date: $
//  $Log: $
//
//
//------------------------------------------------------------------------------


netcdf aot_geo {

//---------
dimensions:
//---------

      Scan = 48;
      Coordinate = 3;
      AlongTrack = 96;
      CrossTrack = 400;


//--------
variables:
//--------


// This is the first array

      ubyte QF1_SCAN_VIIRSAEROGEO(Scan);
            QF1_SCAN_VIIRSAEROGEO:long_name = "Scan-level quality flag";
            QF1_SCAN_VIIRSAEROGEO:units = "none";
            QF1_SCAN_VIIRSAEROGEO:scale_factor = 1.0f;
            QF1_SCAN_VIIRSAEROGEO:add_offset = 0.0f;
            QF1_SCAN_VIIRSAEROGEO:parameter_type = "VIIRS data";
            QF1_SCAN_VIIRSAEROGEO:valid_range = 0ub, 255ub;
            QF1_SCAN_VIIRSAEROGEO:_FillValue = 255ub;

      int64 StartTime(Scan);
            StartTime:long_name = "Start time of scan in IET (1/1/1958)";
            StartTime:units = "microsecond";
            StartTime:scale_factor = 1.0f;
            StartTime:add_offset = 0.0f;
            StartTime:parameter_type = "VIIRS data";
            StartTime:valid_range = 0L, 1000000000000000000L;
            StartTime:_FillValue = -9999L;

      int64 MidTime(Scan);
            MidTime:long_name = "Mid-Time of scan in IET (1/1/1958)";
            MidTime:units = "microsecond";
            MidTime:scale_factor = 1.0f;
            MidTime:add_offset = 0.0f;
            MidTime:parameter_type = "VIIRS data";
            MidTime:valid_range = 0L, 1000000000000000000L;
            MidTime:_FillValue = -9999L;

      float SCPosition(Scan,Coordinate);
            SCPosition:long_name = "Spacecraft position ECR Coordinates";
            SCPosition:units = "meter";
            SCPosition:scale_factor = 1.0f;
            SCPosition:add_offset = 0.0f;
            SCPosition:parameter_type = "VIIRS data";
            SCPosition:valid_range = 0.0f, 1000000.0f;
            SCPosition:_FillValue = -9999.0f;

      float SCVelocity(Scan,Coordinate);
            SCVelocity:long_name = "Spacecraft velocity ECR Coordinates";
            SCVelocity:units = "m/s";
            SCVelocity:scale_factor = 1.0f;
            SCVelocity:add_offset = 0.0f;
            SCVelocity:parameter_type = "VIIRS data";
            SCVelocity:valid_range = 0.0f, 1000000.0f;
            SCVelocity:_FillValue = -9999.0f;

      float SCAttitude(Scan,Coordinate);
            SCAttitude:long_name = "Spacecraft attitude GRF Coordinates";
            SCAttitude:units = "arcsecond";
            SCAttitude:scale_factor = 1.0f;
            SCAttitude:add_offset = 0.0f;
            SCAttitude:parameter_type = "VIIRS data";
            SCAttitude:valid_range = 0.0f, 1000000.0f;
            SCAttitude:_FillValue = -9999.0f;

      float Latitude(AlongTrack,CrossTrack);
            Latitude:long_name = "Latitude of pixel (positive North)";
            Latitude:units = "degree";
            Latitude:scale_factor = 1.0f;
            Latitude:add_offset = 0.0f;
            Latitude:parameter_type = "VIIRS data";
            Latitude:valid_range = -90.0f, 90.0f;
            Latitude:_FillValue = -9999.0f;

      float Longitude(AlongTrack,CrossTrack);
            Longitude:long_name = "Longitude of pixel (positive East)";
            Longitude:units = "degree";
            Longitude:scale_factor = 1.0f;
            Longitude:add_offset = 0.0f;
            Longitude:parameter_type = "VIIRS data";
            Longitude:valid_range = -180.0f, 180.0f;
            Longitude:_FillValue = -9999.0f;

      float SolarZenithAngle(AlongTrack,CrossTrack);
            SolarZenithAngle:long_name = "Zenith angle of sun";
            SolarZenithAngle:units = "degree";
            SolarZenithAngle:scale_factor = 1.0f;
            SolarZenithAngle:add_offset = 0.0f;
            SolarZenithAngle:parameter_type = "VIIRS data";
            SolarZenithAngle:valid_range = 0.0f, 180.0f;
            SolarZenithAngle:_FillValue = -9999.0f;

      float SolarAzimuthAngle(AlongTrack,CrossTrack);
            SolarAzimuthAngle:long_name = "Azimuth angle of sun";
            SolarAzimuthAngle:units = "degree";
            SolarAzimuthAngle:scale_factor = 1.0f;
            SolarAzimuthAngle:add_offset = 0.0f;
            SolarAzimuthAngle:parameter_type = "VIIRS data";
            SolarAzimuthAngle:valid_range = -180.0f, 180.0f;
            SolarAzimuthAngle:_FillValue = -9999.0f;

      float SatelliteZenithAngle(AlongTrack,CrossTrack);
            SatelliteZenithAngle:long_name = "Zenith angle to Satellite";
            SatelliteZenithAngle:units = "degree";
            SatelliteZenithAngle:scale_factor = 1.0f;
            SatelliteZenithAngle:add_offset = 0.0f;
            SatelliteZenithAngle:parameter_type = "VIIRS data";
            SatelliteZenithAngle:valid_range = 0.0f, 70.0f;
            SatelliteZenithAngle:_FillValue = -9999.0f;

      float SatelliteAzimuthAngle(AlongTrack,CrossTrack);
            SatelliteAzimuthAngle:long_name = "Azimuth angle to Satellite";
            SatelliteAzimuthAngle:units = "degree";
            SatelliteAzimuthAngle:scale_factor = 1.0f;
            SatelliteAzimuthAngle:add_offset = 0.0f;
            SatelliteAzimuthAngle:parameter_type = "VIIRS data";
            SatelliteAzimuthAngle:valid_range = -180.0f, 180.0f;
            SatelliteAzimuthAngle:_FillValue = -9999.0f;

      float Height(AlongTrack,CrossTrack);
            Height:long_name = "Ellipsoid-Geoid separation";
            Height:units = "meter";
            Height:scale_factor = 1.0f;
            Height:add_offset = 0.0f;
            Height:parameter_type = "VIIRS data";
            Height:valid_range = 0.0f, 1000000.0f;
            Height:_FillValue = -9999.0f;

      float SatelliteRange(AlongTrack,CrossTrack);
            SatelliteRange:long_name = "Line of sight distance";
            SatelliteRange:units = "meter";
            SatelliteRange:scale_factor = 1.0f;
            SatelliteRange:add_offset = 0.0f;
            SatelliteRange:parameter_type = "VIIRS data";
            SatelliteRange:valid_range = 0.0f, 1000000.0f;
            SatelliteRange:_FillValue = -9999.0f;

// This is the last array

      ubyte QF2_VIIRSAEROGEO(AlongTrack,CrossTrack);
            QF2_VIIRSAEROGEO:long_name = "Pixel-level quality flag";
            QF2_VIIRSAEROGEO:units = "none";
            QF2_VIIRSAEROGEO:scale_factor = 1.0f;
            QF2_VIIRSAEROGEO:add_offset = 0.0f;
            QF2_VIIRSAEROGEO:parameter_type = "VIIRS data";
            QF2_VIIRSAEROGEO:valid_range = 0ub, 255ub;
            QF2_VIIRSAEROGEO:_FillValue = 255ub;


//------------------
// global attributes
//------------------

        :title = "VIIRS MOD GEO granule data file" ;
        :author = "Yi Song IMSG.  Yi.Song@noaa.gov" ;
        :rcsId = "$Id: $" ;


}
